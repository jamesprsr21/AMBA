Protocol are nothing but set of rules by which we can communicate between master and slave.
There are two types of Protocol. 1> Onchip protocol ; 2>Offchip/Peripheral Protocol.
The SoC has several functional blocks that use AMBA protocols like AXI4 and AXI3 to communicate with each other.

AMBA stands for Advanced Microcontroller Bus Architecture
  It is a onchip protocol. Which is used to connect functional blocks which are on the chip(SOC).
Essentially, AMBA protocols define how functional blocks communicate with each other.
