AXI stands for Advanced eXtensible Interface.
  It is a high-performance, parallel bus that connects processor cores to on-chip peripheral circuits.
  A high-performance, point-to-point, master-slave parallel bus that connects processor cores to on-chip peripheral circuits
